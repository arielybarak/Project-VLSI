/*------------------------------------------------------------------------------
 * File          : one_hot_encoder.sv
 * Project       : RTL
 * Author        : epabab
 * Creation date : Sep 18, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

module one_hot_encoder #() ();

endmodule